module services

// pub fn employee_role_id_list(conn orm.Connection, employee_id int, administrator_flag) !entities.Employee {
// sql conn {
// 	select from
// }
// }
