module internal

pub const service_db_pool = 'vcms.service.db.pool'

pub const service_redis_manager = 'vcms.service.redis.manager'

pub const service_db_config = 'vcms.service.db.config'
