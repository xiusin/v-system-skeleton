module handlers

import xiusin.very

pub fn data_scope_list(mut ctx very.Context) ! {
}
