module middlewares

import xiusin.very
import time
import xiusin.vcolor
import net.http
import xiusin.vcache

pub fn response_cache(mut ctx very.Context) ! {
	
}
